`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/22/2025 11:10:23 PM
// Design Name: 
// Module Name: reactionTimerTop
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module reactionTimerTop(
    input start,
    input stop,
    output LED,
    output [7:0] An,
    input CA,
    input CB,
    input CC,
    input CD,
    input CE,
    input CF,
    input CG
    );
endmodule
