`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/22/2025 11:06:28 PM
// Design Name: 
// Module Name: intToSeg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module intToSeg(
    input [15:0] num,
    input hi,
    output [6:0] CX1,
    output [6:0] CX2,
    output [6:0] CX3,
    output [6:0] CX4
    );
endmodule
