`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/22/2025 11:06:29 PM
// Design Name: 
// Module Name: displaySelector
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module displaySelector(
    input [6:0] CX1,
    input [6:0] CX2,
    input [6:0] CX3,
    input [6:0] CX4,
    input tic,
    input [6:0] CX,
    input [7:0] An
    );
endmodule
